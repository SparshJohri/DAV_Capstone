module FullFFT #(SAMPLES = 8, WIDTH = 16)
(
	input [WIDTH-1:0] inputs [SAMPLES-1:0],
	input clk,
	output [WIDTH-1:0] outputs [SAMPLES-1:0]
);

	logic [WIDTH-1:0] newRow [SAMPLES-1:0];


endmodule
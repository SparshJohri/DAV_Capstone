module vga_top_tb
(
	
);



endmodule
module Ping_Pong_RAM
(

);


/*

*/



endmodule
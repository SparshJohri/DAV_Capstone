module twiddleFactorCalculator #(parameter SAMPLES=8, WIDTH = 8)
(
	input [$clog2(SAMPLES)-1:0] which_factor,
	output [(WIDTH-1):0] result
);

		logic [(WIDTH/2)-1:0] result_real;
		logic [(WIDTH/2)-1:0] result_imag;
		
		
		logic [(WIDTH/2)-1:0] lookupTableCosines [127:0];
		logic [(WIDTH/2)-1:0] lookupTableSines   [127:0];
		
		int x;
		
		assign x = (256>>($clog2(SAMPLES)))*(which_factor);
		
		assign result_real = lookupTableCosines[(which_factor)*(256>>($clog2(SAMPLES)))];
		assign result_imag = lookupTableSines[(which_factor)*(256>>($clog2(SAMPLES)))];
		
		assign result[(WIDTH-1):(WIDTH/2)] = result_imag;
		assign result[((WIDTH/2) -1):0] = result_real;
		
		
		
		initial
		begin
			lookupTableCosines[0] = (2**( (WIDTH/2) -1))*1.0;
			lookupTableCosines[1] = (2**( (WIDTH/2) -1))*0.999;
			lookupTableCosines[2] = (2**( (WIDTH/2) -1))*0.998;
			lookupTableCosines[3] = (2**( (WIDTH/2) -1))*0.997;
			lookupTableCosines[4] = (2**( (WIDTH/2) -1))*0.995;
			lookupTableCosines[5] = (2**( (WIDTH/2) -1))*0.992;
			lookupTableCosines[6] = (2**( (WIDTH/2) -1))*0.989;
			lookupTableCosines[7] = (2**( (WIDTH/2) -1))*0.985;
			lookupTableCosines[8] = (2**( (WIDTH/2) -1))*0.98;
			lookupTableCosines[9] = (2**( (WIDTH/2) -1))*0.975;
			lookupTableCosines[10] = (2**( (WIDTH/2) -1))*0.97;
			lookupTableCosines[11] = (2**( (WIDTH/2) -1))*0.963;
			lookupTableCosines[12] = (2**( (WIDTH/2) -1))*0.956;
			lookupTableCosines[13] = (2**( (WIDTH/2) -1))*0.949;
			lookupTableCosines[14] = (2**( (WIDTH/2) -1))*0.941;
			lookupTableCosines[15] = (2**( (WIDTH/2) -1))*0.932;
			lookupTableCosines[16] = (2**( (WIDTH/2) -1))*0.923;
			lookupTableCosines[17] = (2**( (WIDTH/2) -1))*0.914;
			lookupTableCosines[18] = (2**( (WIDTH/2) -1))*0.903;
			lookupTableCosines[19] = (2**( (WIDTH/2) -1))*0.893;
			lookupTableCosines[20] = (2**( (WIDTH/2) -1))*0.881;
			lookupTableCosines[21] = (2**( (WIDTH/2) -1))*0.87;
			lookupTableCosines[22] = (2**( (WIDTH/2) -1))*0.857;
			lookupTableCosines[23] = (2**( (WIDTH/2) -1))*0.844;
			lookupTableCosines[24] = (2**( (WIDTH/2) -1))*0.831;
			lookupTableCosines[25] = (2**( (WIDTH/2) -1))*0.817;
			lookupTableCosines[26] = (2**( (WIDTH/2) -1))*0.803;
			lookupTableCosines[27] = (2**( (WIDTH/2) -1))*0.788;
			lookupTableCosines[28] = (2**( (WIDTH/2) -1))*0.773;
			lookupTableCosines[29] = (2**( (WIDTH/2) -1))*0.757;
			lookupTableCosines[30] = (2**( (WIDTH/2) -1))*0.74;
			lookupTableCosines[31] = (2**( (WIDTH/2) -1))*0.724;
			lookupTableCosines[32] = (2**( (WIDTH/2) -1))*0.707;
			lookupTableCosines[33] = (2**( (WIDTH/2) -1))*0.689;
			lookupTableCosines[34] = (2**( (WIDTH/2) -1))*0.671;
			lookupTableCosines[35] = (2**( (WIDTH/2) -1))*0.653;
			lookupTableCosines[36] = (2**( (WIDTH/2) -1))*0.634;
			lookupTableCosines[37] = (2**( (WIDTH/2) -1))*0.615;
			lookupTableCosines[38] = (2**( (WIDTH/2) -1))*0.595;
			lookupTableCosines[39] = (2**( (WIDTH/2) -1))*0.575;
			lookupTableCosines[40] = (2**( (WIDTH/2) -1))*0.555;
			lookupTableCosines[41] = (2**( (WIDTH/2) -1))*0.534;
			lookupTableCosines[42] = (2**( (WIDTH/2) -1))*0.514;
			lookupTableCosines[43] = (2**( (WIDTH/2) -1))*0.492;
			lookupTableCosines[44] = (2**( (WIDTH/2) -1))*0.471;
			lookupTableCosines[45] = (2**( (WIDTH/2) -1))*0.449;
			lookupTableCosines[46] = (2**( (WIDTH/2) -1))*0.427;
			lookupTableCosines[47] = (2**( (WIDTH/2) -1))*0.405;
			lookupTableCosines[48] = (2**( (WIDTH/2) -1))*0.382;
			lookupTableCosines[49] = (2**( (WIDTH/2) -1))*0.359;
			lookupTableCosines[50] = (2**( (WIDTH/2) -1))*0.336;
			lookupTableCosines[51] = (2**( (WIDTH/2) -1))*0.313;
			lookupTableCosines[52] = (2**( (WIDTH/2) -1))*0.29;
			lookupTableCosines[53] = (2**( (WIDTH/2) -1))*0.266;
			lookupTableCosines[54] = (2**( (WIDTH/2) -1))*0.242;
			lookupTableCosines[55] = (2**( (WIDTH/2) -1))*0.219;
			lookupTableCosines[56] = (2**( (WIDTH/2) -1))*0.195;
			lookupTableCosines[57] = (2**( (WIDTH/2) -1))*0.17;
			lookupTableCosines[58] = (2**( (WIDTH/2) -1))*0.146;
			lookupTableCosines[59] = (2**( (WIDTH/2) -1))*0.122;
			lookupTableCosines[60] = (2**( (WIDTH/2) -1))*0.098;
			lookupTableCosines[61] = (2**( (WIDTH/2) -1))*0.073;
			lookupTableCosines[62] = (2**( (WIDTH/2) -1))*0.049;
			lookupTableCosines[63] = (2**( (WIDTH/2) -1))*0.024;
			lookupTableCosines[64] = (2**( (WIDTH/2) -1))*0.0;
			lookupTableCosines[65] = (2**( (WIDTH/2) -1))*-0.024;
			lookupTableCosines[66] = (2**( (WIDTH/2) -1))*-0.049;
			lookupTableCosines[67] = (2**( (WIDTH/2) -1))*-0.073;
			lookupTableCosines[68] = (2**( (WIDTH/2) -1))*-0.098;
			lookupTableCosines[69] = (2**( (WIDTH/2) -1))*-0.122;
			lookupTableCosines[70] = (2**( (WIDTH/2) -1))*-0.146;
			lookupTableCosines[71] = (2**( (WIDTH/2) -1))*-0.17;
			lookupTableCosines[72] = (2**( (WIDTH/2) -1))*-0.195;
			lookupTableCosines[73] = (2**( (WIDTH/2) -1))*-0.219;
			lookupTableCosines[74] = (2**( (WIDTH/2) -1))*-0.242;
			lookupTableCosines[75] = (2**( (WIDTH/2) -1))*-0.266;
			lookupTableCosines[76] = (2**( (WIDTH/2) -1))*-0.29;
			lookupTableCosines[77] = (2**( (WIDTH/2) -1))*-0.313;
			lookupTableCosines[78] = (2**( (WIDTH/2) -1))*-0.336;
			lookupTableCosines[79] = (2**( (WIDTH/2) -1))*-0.359;
			lookupTableCosines[80] = (2**( (WIDTH/2) -1))*-0.382;
			lookupTableCosines[81] = (2**( (WIDTH/2) -1))*-0.405;
			lookupTableCosines[82] = (2**( (WIDTH/2) -1))*-0.427;
			lookupTableCosines[83] = (2**( (WIDTH/2) -1))*-0.449;
			lookupTableCosines[84] = (2**( (WIDTH/2) -1))*-0.471;
			lookupTableCosines[85] = (2**( (WIDTH/2) -1))*-0.492;
			lookupTableCosines[86] = (2**( (WIDTH/2) -1))*-0.514;
			lookupTableCosines[87] = (2**( (WIDTH/2) -1))*-0.534;
			lookupTableCosines[88] = (2**( (WIDTH/2) -1))*-0.555;
			lookupTableCosines[89] = (2**( (WIDTH/2) -1))*-0.575;
			lookupTableCosines[90] = (2**( (WIDTH/2) -1))*-0.595;
			lookupTableCosines[91] = (2**( (WIDTH/2) -1))*-0.615;
			lookupTableCosines[92] = (2**( (WIDTH/2) -1))*-0.634;
			lookupTableCosines[93] = (2**( (WIDTH/2) -1))*-0.653;
			lookupTableCosines[94] = (2**( (WIDTH/2) -1))*-0.671;
			lookupTableCosines[95] = (2**( (WIDTH/2) -1))*-0.689;
			lookupTableCosines[96] = (2**( (WIDTH/2) -1))*-0.707;
			lookupTableCosines[97] = (2**( (WIDTH/2) -1))*-0.724;
			lookupTableCosines[98] = (2**( (WIDTH/2) -1))*-0.74;
			lookupTableCosines[99] = (2**( (WIDTH/2) -1))*-0.757;
			lookupTableCosines[100] = (2**( (WIDTH/2) -1))*-0.773;
			lookupTableCosines[101] = (2**( (WIDTH/2) -1))*-0.788;
			lookupTableCosines[102] = (2**( (WIDTH/2) -1))*-0.803;
			lookupTableCosines[103] = (2**( (WIDTH/2) -1))*-0.817;
			lookupTableCosines[104] = (2**( (WIDTH/2) -1))*-0.831;
			lookupTableCosines[105] = (2**( (WIDTH/2) -1))*-0.844;
			lookupTableCosines[106] = (2**( (WIDTH/2) -1))*-0.857;
			lookupTableCosines[107] = (2**( (WIDTH/2) -1))*-0.87;
			lookupTableCosines[108] = (2**( (WIDTH/2) -1))*-0.881;
			lookupTableCosines[109] = (2**( (WIDTH/2) -1))*-0.893;
			lookupTableCosines[110] = (2**( (WIDTH/2) -1))*-0.903;
			lookupTableCosines[111] = (2**( (WIDTH/2) -1))*-0.914;
			lookupTableCosines[112] = (2**( (WIDTH/2) -1))*-0.923;
			lookupTableCosines[113] = (2**( (WIDTH/2) -1))*-0.932;
			lookupTableCosines[114] = (2**( (WIDTH/2) -1))*-0.941;
			lookupTableCosines[115] = (2**( (WIDTH/2) -1))*-0.949;
			lookupTableCosines[116] = (2**( (WIDTH/2) -1))*-0.956;
			lookupTableCosines[117] = (2**( (WIDTH/2) -1))*-0.963;
			lookupTableCosines[118] = (2**( (WIDTH/2) -1))*-0.97;
			lookupTableCosines[119] = (2**( (WIDTH/2) -1))*-0.975;
			lookupTableCosines[120] = (2**( (WIDTH/2) -1))*-0.98;
			lookupTableCosines[121] = (2**( (WIDTH/2) -1))*-0.985;
			lookupTableCosines[122] = (2**( (WIDTH/2) -1))*-0.989;
			lookupTableCosines[123] = (2**( (WIDTH/2) -1))*-0.992;
			lookupTableCosines[124] = (2**( (WIDTH/2) -1))*-0.995;
			lookupTableCosines[125] = (2**( (WIDTH/2) -1))*-0.997;
			lookupTableCosines[126] = (2**( (WIDTH/2) -1))*-0.998;
			lookupTableCosines[127] = (2**( (WIDTH/2) -1))*-0.999;

			lookupTableSines[0] = (2**( (WIDTH/2) -1))*0.0;
			lookupTableSines[1] = (2**( (WIDTH/2) -1))*0.024;
			lookupTableSines[2] = (2**( (WIDTH/2) -1))*0.049;
			lookupTableSines[3] = (2**( (WIDTH/2) -1))*0.073;
			lookupTableSines[4] = (2**( (WIDTH/2) -1))*0.098;
			lookupTableSines[5] = (2**( (WIDTH/2) -1))*0.122;
			lookupTableSines[6] = (2**( (WIDTH/2) -1))*0.146;
			lookupTableSines[7] = (2**( (WIDTH/2) -1))*0.17;
			lookupTableSines[8] = (2**( (WIDTH/2) -1))*0.195;
			lookupTableSines[9] = (2**( (WIDTH/2) -1))*0.219;
			lookupTableSines[10] = (2**( (WIDTH/2) -1))*0.242;
			lookupTableSines[11] = (2**( (WIDTH/2) -1))*0.266;
			lookupTableSines[12] = (2**( (WIDTH/2) -1))*0.29;
			lookupTableSines[13] = (2**( (WIDTH/2) -1))*0.313;
			lookupTableSines[14] = (2**( (WIDTH/2) -1))*0.336;
			lookupTableSines[15] = (2**( (WIDTH/2) -1))*0.359;
			lookupTableSines[16] = (2**( (WIDTH/2) -1))*0.382;
			lookupTableSines[17] = (2**( (WIDTH/2) -1))*0.405;
			lookupTableSines[18] = (2**( (WIDTH/2) -1))*0.427;
			lookupTableSines[19] = (2**( (WIDTH/2) -1))*0.449;
			lookupTableSines[20] = (2**( (WIDTH/2) -1))*0.471;
			lookupTableSines[21] = (2**( (WIDTH/2) -1))*0.492;
			lookupTableSines[22] = (2**( (WIDTH/2) -1))*0.514;
			lookupTableSines[23] = (2**( (WIDTH/2) -1))*0.534;
			lookupTableSines[24] = (2**( (WIDTH/2) -1))*0.555;
			lookupTableSines[25] = (2**( (WIDTH/2) -1))*0.575;
			lookupTableSines[26] = (2**( (WIDTH/2) -1))*0.595;
			lookupTableSines[27] = (2**( (WIDTH/2) -1))*0.615;
			lookupTableSines[28] = (2**( (WIDTH/2) -1))*0.634;
			lookupTableSines[29] = (2**( (WIDTH/2) -1))*0.653;
			lookupTableSines[30] = (2**( (WIDTH/2) -1))*0.671;
			lookupTableSines[31] = (2**( (WIDTH/2) -1))*0.689;
			lookupTableSines[32] = (2**( (WIDTH/2) -1))*0.707;
			lookupTableSines[33] = (2**( (WIDTH/2) -1))*0.724;
			lookupTableSines[34] = (2**( (WIDTH/2) -1))*0.74;
			lookupTableSines[35] = (2**( (WIDTH/2) -1))*0.757;
			lookupTableSines[36] = (2**( (WIDTH/2) -1))*0.773;
			lookupTableSines[37] = (2**( (WIDTH/2) -1))*0.788;
			lookupTableSines[38] = (2**( (WIDTH/2) -1))*0.803;
			lookupTableSines[39] = (2**( (WIDTH/2) -1))*0.817;
			lookupTableSines[40] = (2**( (WIDTH/2) -1))*0.831;
			lookupTableSines[41] = (2**( (WIDTH/2) -1))*0.844;
			lookupTableSines[42] = (2**( (WIDTH/2) -1))*0.857;
			lookupTableSines[43] = (2**( (WIDTH/2) -1))*0.87;
			lookupTableSines[44] = (2**( (WIDTH/2) -1))*0.881;
			lookupTableSines[45] = (2**( (WIDTH/2) -1))*0.893;
			lookupTableSines[46] = (2**( (WIDTH/2) -1))*0.903;
			lookupTableSines[47] = (2**( (WIDTH/2) -1))*0.914;
			lookupTableSines[48] = (2**( (WIDTH/2) -1))*0.923;
			lookupTableSines[49] = (2**( (WIDTH/2) -1))*0.932;
			lookupTableSines[50] = (2**( (WIDTH/2) -1))*0.941;
			lookupTableSines[51] = (2**( (WIDTH/2) -1))*0.949;
			lookupTableSines[52] = (2**( (WIDTH/2) -1))*0.956;
			lookupTableSines[53] = (2**( (WIDTH/2) -1))*0.963;
			lookupTableSines[54] = (2**( (WIDTH/2) -1))*0.97;
			lookupTableSines[55] = (2**( (WIDTH/2) -1))*0.975;
			lookupTableSines[56] = (2**( (WIDTH/2) -1))*0.98;
			lookupTableSines[57] = (2**( (WIDTH/2) -1))*0.985;
			lookupTableSines[58] = (2**( (WIDTH/2) -1))*0.989;
			lookupTableSines[59] = (2**( (WIDTH/2) -1))*0.992;
			lookupTableSines[60] = (2**( (WIDTH/2) -1))*0.995;
			lookupTableSines[61] = (2**( (WIDTH/2) -1))*0.997;
			lookupTableSines[62] = (2**( (WIDTH/2) -1))*0.998;
			lookupTableSines[63] = (2**( (WIDTH/2) -1))*0.999;
			lookupTableSines[64] = (2**( (WIDTH/2) -1))*1.0;
			lookupTableSines[65] = (2**( (WIDTH/2) -1))*0.999;
			lookupTableSines[66] = (2**( (WIDTH/2) -1))*0.998;
			lookupTableSines[67] = (2**( (WIDTH/2) -1))*0.997;
			lookupTableSines[68] = (2**( (WIDTH/2) -1))*0.995;
			lookupTableSines[69] = (2**( (WIDTH/2) -1))*0.992;
			lookupTableSines[70] = (2**( (WIDTH/2) -1))*0.989;
			lookupTableSines[71] = (2**( (WIDTH/2) -1))*0.985;
			lookupTableSines[72] = (2**( (WIDTH/2) -1))*0.98;
			lookupTableSines[73] = (2**( (WIDTH/2) -1))*0.975;
			lookupTableSines[74] = (2**( (WIDTH/2) -1))*0.97;
			lookupTableSines[75] = (2**( (WIDTH/2) -1))*0.963;
			lookupTableSines[76] = (2**( (WIDTH/2) -1))*0.956;
			lookupTableSines[77] = (2**( (WIDTH/2) -1))*0.949;
			lookupTableSines[78] = (2**( (WIDTH/2) -1))*0.941;
			lookupTableSines[79] = (2**( (WIDTH/2) -1))*0.932;
			lookupTableSines[80] = (2**( (WIDTH/2) -1))*0.923;
			lookupTableSines[81] = (2**( (WIDTH/2) -1))*0.914;
			lookupTableSines[82] = (2**( (WIDTH/2) -1))*0.903;
			lookupTableSines[83] = (2**( (WIDTH/2) -1))*0.893;
			lookupTableSines[84] = (2**( (WIDTH/2) -1))*0.881;
			lookupTableSines[85] = (2**( (WIDTH/2) -1))*0.87;
			lookupTableSines[86] = (2**( (WIDTH/2) -1))*0.857;
			lookupTableSines[87] = (2**( (WIDTH/2) -1))*0.844;
			lookupTableSines[88] = (2**( (WIDTH/2) -1))*0.831;
			lookupTableSines[89] = (2**( (WIDTH/2) -1))*0.817;
			lookupTableSines[90] = (2**( (WIDTH/2) -1))*0.803;
			lookupTableSines[91] = (2**( (WIDTH/2) -1))*0.788;
			lookupTableSines[92] = (2**( (WIDTH/2) -1))*0.773;
			lookupTableSines[93] = (2**( (WIDTH/2) -1))*0.757;
			lookupTableSines[94] = (2**( (WIDTH/2) -1))*0.74;
			lookupTableSines[95] = (2**( (WIDTH/2) -1))*0.724;
			lookupTableSines[96] = (2**( (WIDTH/2) -1))*0.707;
			lookupTableSines[97] = (2**( (WIDTH/2) -1))*0.689;
			lookupTableSines[98] = (2**( (WIDTH/2) -1))*0.671;
			lookupTableSines[99] = (2**( (WIDTH/2) -1))*0.653;
			lookupTableSines[100] = (2**( (WIDTH/2) -1))*0.634;
			lookupTableSines[101] = (2**( (WIDTH/2) -1))*0.615;
			lookupTableSines[102] = (2**( (WIDTH/2) -1))*0.595;
			lookupTableSines[103] = (2**( (WIDTH/2) -1))*0.575;
			lookupTableSines[104] = (2**( (WIDTH/2) -1))*0.555;
			lookupTableSines[105] = (2**( (WIDTH/2) -1))*0.534;
			lookupTableSines[106] = (2**( (WIDTH/2) -1))*0.514;
			lookupTableSines[107] = (2**( (WIDTH/2) -1))*0.492;
			lookupTableSines[108] = (2**( (WIDTH/2) -1))*0.471;
			lookupTableSines[109] = (2**( (WIDTH/2) -1))*0.449;
			lookupTableSines[110] = (2**( (WIDTH/2) -1))*0.427;
			lookupTableSines[111] = (2**( (WIDTH/2) -1))*0.405;
			lookupTableSines[112] = (2**( (WIDTH/2) -1))*0.382;
			lookupTableSines[113] = (2**( (WIDTH/2) -1))*0.359;
			lookupTableSines[114] = (2**( (WIDTH/2) -1))*0.336;
			lookupTableSines[115] = (2**( (WIDTH/2) -1))*0.313;
			lookupTableSines[116] = (2**( (WIDTH/2) -1))*0.29;
			lookupTableSines[117] = (2**( (WIDTH/2) -1))*0.266;
			lookupTableSines[118] = (2**( (WIDTH/2) -1))*0.242;
			lookupTableSines[119] = (2**( (WIDTH/2) -1))*0.219;
			lookupTableSines[120] = (2**( (WIDTH/2) -1))*0.195;
			lookupTableSines[121] = (2**( (WIDTH/2) -1))*0.17;
			lookupTableSines[122] = (2**( (WIDTH/2) -1))*0.146;
			lookupTableSines[123] = (2**( (WIDTH/2) -1))*0.122;
			lookupTableSines[124] = (2**( (WIDTH/2) -1))*0.098;
			lookupTableSines[125] = (2**( (WIDTH/2) -1))*0.073;
			lookupTableSines[126] = (2**( (WIDTH/2) -1))*0.049;
			lookupTableSines[127] = (2**( (WIDTH/2) -1))*0.024;		
	end

endmodule
module Microphone_testing
(

);



endmodule